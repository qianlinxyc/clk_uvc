package clk_uvc_pkg;
    import uvm_pkg::*;

    `include "clk_uvc_cfg.sv"
    `include "clk_uvc_drv.sv"
    `include "clk_uvc_agt.sv"
endpackage : clk_uvc_pkg
